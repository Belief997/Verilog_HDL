
module  FretoFre(  
    input                                   clk,  
    input                                   rst_n,  
  
    output                                  clk_2M//,  
//    output      reg         [4:0]               Count  
);  
  
//??????????????????????????????????????????????????????????????????-????????????????  
//              ???????  
reg           [4:0]               Count; 
initial Count = 'b0; 
always @ (posedge clk or negedge rst_n)           
begin  
    if(!rst_n)  
        Count <= 'd0;  
    else if(Count >= 5'd24)  
        Count <= 'd0;  
    else  
        Count <= Count + 1'b1;  
end  
  
//???????????????????????????????????????????????????????????????????????????????????  
//  ??????????????12/25??????  
reg                             Pos_clk;  
always @ (posedge clk or negedge rst_n)  
begin  
    if(!rst_n)  
        Pos_clk <= 'd0;  
    else if(Count >= 5'd13)  
        Pos_clk <= 1'b1;  
    else  
        Pos_clk <= 'd0;  
end  

//???????????????????????????????????????????????????????????????????????????????????  
//??????????????12/25??????  
reg                             Neg_clk;  
always @ (negedge clk or negedge rst_n)  
begin  
    if(!rst_n)  
        Neg_clk <= 'd0;  
    else if(Count >= 5'd13)  
        Neg_clk <= 1'b1;  
    else  
        Neg_clk <= 'd0;  
end  
  
//???????????????????????????????????????????????????????????????????????????????????  
//          ???  
assign  clk_2M = Pos_clk | Neg_clk;  
  
endmodule 