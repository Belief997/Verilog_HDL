`timescale 1ns/1ps
module tb;
    	reg clk;
//	wire signed [7:0] Out;
	reg key1, key2 ,key3, key4, key5, key6, key7, key0;
	reg signed [11:0] m ;
	wire pwm;
/*	wire signed [7:0] data = 8'hc0;
	wire pwmp, pwmn;*/
//    reg [23:0] freq;
//    wire [23:0] phaseShift = 24'b0;
//    wire clkEn = 1'b1;
//    wire signed [11:0] out;
//    initial begin
//        clk = 1'b1;
//        freq = 24'd1678;
//        /*#10010 freq = 24'h08_0000;
//        #20000 freq = 24'h0C_0000;
//        #30000 freq = 24'h10_0000;
//        #40000 freq = 24'h18_0000;
//        #50000 freq = 24'h20_0000;
//        #60000 freq = 24'h30_0000;*/
//        //#70000 $stop();
//    end
//    always begin
//        #5 clk = ~clk;
//    end    
//    dds #( 
//	.PHASE_W (24), 
//	.DATA_W (12), 
//	.TABLE_AW  (12),
//	.MEM_FILE  ("SineTable12X12.dat")
//) dds_inst (
//       .FreqWord(freq),
//       .PhaseShift(phaseShift),
//       .clk(clk),
//       .ClkEn(clkEn),
//       .Out(out)) ;

initial begin 
	clk = 1'b0;
	key1= 1'b0;
	key2 =1'b0;
	key3= 1'b0;
	key4= 1'b0;
	key5= 1'b0;
	key6= 1'b0;
	key7= 1'b0;
	key0 = 1'b0;
	m = 12'sd1024;//(0.5) //1844(0.9);//2048(-1);
end
always begin
	#999999  key1 = 1'b1;
	#50 key1 = 1'b0;
	#99  key1 = 1'b1;
	#50 key1 = 1'b0;
	#999  key1 = 1'b1;
	#50 key1 = 1'b0;
	#999  key1 = 1'b1;
	#50 key1 = 1'b0;
	#99  key1 = 1'b1;
	#50 key1 = 1'b0;
	//#50 m = m - 12'sd204;
end
always begin 
	#5 clk =~clk;
end

always begin
	#999999  key7 = 1'b1;
	#50 key7 = 1'b0;
	#99  key7 = 1'b1;
	#50 key7 = 1'b0;
	#999  key7 = 1'b1;
	#50 key7 = 1'b0;
	#999  key7 = 1'b1;
	#50 key7 = 1'b0;
	#99  key7 = 1'b1;
	#50 key7 = 1'b0;
end
//PWM the_pwm( 
//	.clk(clk), .rst(1'b0), 
//	.data(data), 
//	.pwm(pwm)
//);



top the_top(
	.clk(clk),
	.rst(1'b0),
	.m0(m),
	.key1(key1), .key2(key2) ,.key3(key3), .key4(key4), .key5(key5), .key6(key6), .key7(key7), .key0(key0),
	.pwm(pwm)
	);
endmodule

	