//10kbps
//module LFSR(
//	input clk, en,
//	output reg out
//);
//initial out = 'b0;
//always@(posedge clk)begin
//	if(en) out <= ~out;
//
//end
//
//
//
//
//
//endmodule 
//
//

//W is the highest pow 
//MASK :  its LSB is not cared 
module LFSR#( parameter W = 8, parameter [W:0] MASK = 32'h11c //, parameter WO = W
)(
	input clk, clken,
	output reg [W - 1 : 0] lfsr
);
	initial lfsr = 'b1;

	always@(posedge clk)begin
		if(clken)begin
			if(lfsr[0]) lfsr <= (lfsr >> 1) ^ (MASK >> 1);
			else lfsr <= (lfsr >> 1);
		end
	end
endmodule 
