
module my_iir(
	input clk,
	input signed [31:0] in,
	output signed [31:0] out

);
	wire signed [31:0] y1x2_1, y2x3_1, y3x4_1,y4x5_1, out_1;
	wire signed [31:0] y1x2_2, y2x3_2, y3x4_2,y4x5_2, out_2;
	wire signed [31:0] y1x2_3, y2x3_3, y3x4_3,y4x5_3, out_3;
	wire signed [31:0] y1x2_4, y2x3_4, y3x4_4,y4x5_4, out_4;
	wire signed [31:0] y1x2_5;
//	reg signed [31:0] sec12, sec23, sec34, sec45, sec56;
	/*(* mark_debug = "true" *)*/reg signed [31:0] the_in;
	
	reg [3:0] cnten;
initial begin cnten = 4'b1; the_in = 'b0; /*sec12 ='b0;sec23 ='b0;sec34 ='b0;sec45 ='b0;sec56 ='b0; */end
always @(posedge clk) begin
	if((cnten!=4'd10))
		cnten <= cnten + 1'b1;
	else if (cnten == 4'd10) begin
		cnten <= 4'd10;
	end 
end

always @(posedge clk) begin
    the_in <= in;
//    sec12 <= y1x2;
//    sec23 <= y2x3;
//    sec34 <= y3x4;
//    sec45 <= y4x5;
////    sec56 <= y5x6;
end
//assi

wire en=(cnten == 4'd10);



//////Fs 4 Order 44 Sec22 Butter
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0063346527219021107     ),
	.B1(2        *0.0063346527219021107     ),
	.B2(1*0.0063346527219021107     ),
	.A1(-1.9633665835404945       ),
	.A2( 0.98870519442810278      )
) p1sec1 (
	.clk(clk),.en(en),
	.in(the_in),
	.out(y1x2_1)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.006264081407241791      ),
	.B1(2*0.006264081407241791      ),
	.B2(1*0.006264081407241791      ),
	.A1(-1.9414936621597327       ),
	.A2( 0.96654998778869983      )
) p1sec2 (
	.clk(clk),.en(en),
	.in(y1x2_1),
	.out(y2x3_1)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.006195587382611294      ),
	.B1(2*0.006195587382611294      ),
	.B2(1*0.006195587382611294      ),
	.A1(-1.9202645774670937       ),
	.A2( 0.94504692699753901      )
) p1sec3 (
	.clk(clk),.en(en),
	.in(y2x3_1),
	.out(y3x4_1)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0061294239634460557     ),
	.B1(2*0.0061294239634460557     ),
	.B2(1*0.0061294239634460557     ),
	.A1(-1.8997578422213444       ),
	.A2( 0.92427553807512852      )    
) p1sec4(
	.clk(clk),.en(en),
	.in(y3x4_1),
	.out(y4x5_1)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0060658167028956218     ),
	.B1(2*0.0060658167028956218     ),
	.B2(1*0.0060658167028956218     ),
	.A1(-1.8800433645194357       ),
	.A2( 0.90430663133101807      )    
) p1sec5(
	.clk(clk),.en(en),
	.in(y4x5_1),
	.out(out_1)
);
///// part1 end
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0060049651021757263     ),
	.B1(2*0.0060049651021757263     ),
	.B2(1*0.0060049651021757263     ),
	.A1(-1.8611829779041897       ),
	.A2( 0.8852028383128927       )
) p2sec1 (
	.clk(clk),.en(en),
	.in(out_1),
	.out(y1x2_2)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0059470444625051248     ),
	.B1(2*0.0059470444625051248     ),
	.B2(1*0.0059470444625051248     ),
	.A1(-1.8432310153548674        ),
	.A2( 0.86701919320488796      )
) p2sec2 (
	.clk(clk),.en(en),
	.in(y1x2_2),
	.out(y2x3_2)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0058922078155218636     ),
	.B1(2*0.0058922078155218636     ),
	.B2(1*0.0058922078155218636     ),
	.A1(-1.8262349076017006       ),
	.A2( 0.84980373886378802      )
) p2sec3 (
	.clk(clk),.en(en),
	.in(y2x3_2),
	.out(y3x4_2)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.005840587878771019      ),
	.B1(2*0.005840587878771019      ),
	.B2(1*0.005840587878771019      ),
	.A1(-1.8102357892110954       ),
	.A2( 0.83359814072617955      )    
) p2sec4(
	.clk(clk),.en(en),
	.in(y3x4_2),
	.out(y4x5_2)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0057922989920710403     ),
	.B1(2*0.0057922989920710403     ),
	.B2(1*0.0057922989920710403     ),
	.A1(-1.7952690987443376       ),
	.A2( 0.81843829471262197      )    
) p2sec5(
	.clk(clk),.en(en),
	.in(y4x5_2),
	.out(out_2)
);
//part 2 end
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0057474389990412322     ),
	.B1(2*0.0057474389990412322     ),
	.B2(1*0.0057474389990412322     ),
	.A1(-1.7813651619195046       ),
	.A2( 0.8043549179156696       )
) p3sec1 (
	.clk(clk),.en(en),
	.in(out_2),
	.out(y1x2_3)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0057060910456511217     ),
	.B1(2 *0.0057060910456511217     ),
	.B2(1*0.0057060910456511217     ),
	.A1(-1.768549749055079         ),
	.A2( 0.79137411323768347      )
) p3sec2 (
	.clk(clk),.en(en),
	.in(y1x2_3),
	.out(y2x3_3)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0056683252742563642     ),
	.B1(2*0.0056683252742563642     ),
	.B2(1*0.0056683252742563642     ),
	.A1(-1.7568446001205955       ),
	.A2( 0.77951790121762088      )
) p3sec3 (
	.clk(clk),.en(en),
	.in(y2x3_3),
	.out(y3x4_3)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0056342003972003939     ),
	.B1(2*0.0056342003972003939     ),
	.B2(1*0.0056342003972003939     ),
	.A1(-1.7462679124598073       ),
	.A2( 0.76880471404860895      )    
) p3sec4(
	.clk(clk),.en(en),
	.in(y3x4_3),
	.out(y4x5_3)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0056037651387159416     ),
	.B1(2*0.0056037651387159416     ),
	.B2(1*0.0056037651387159416     ),
	.A1(-1.7368347876946271       ),
	.A2( 0.75924984824949082      )    
) p3sec5(
	.clk(clk),.en(en),
	.in(y4x5_3),
	.out(out_3)
);
//part 3 end
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.00557705953761721       ),
	.B1(2*0.00557705953761721       ),
	.B2(1*0.00557705953761721       ),
	.A1(-1.7285576354824268       ),
	.A2( 0.7508658736328957       )
) p4sec1 (
	.clk(clk),.en(en),
	.in(out_3),
	.out(y1x2_4)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0055541161062122668     ),
	.B1(2*0.0055541161062122668     ),
	.B2(1*0.0055541161062122668     ),
	.A1(-1.7214465327101358       ),
	.A2( 0.74366299713498485      )
) p4sec2 (
	.clk(clk),.en(en),
	.in(y1x2_4),
	.out(y2x3_4)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0055349608430775212     ),
	.B1(2*0.0055349608430775212     ),
	.B2(1*0.0055349608430775212     ),
	.A1(-1.7155095373942519       ),
	.A2( 0.73764938076656184      )
) p4sec3 (
	.clk(clk),.en(en),
	.in(y2x3_4),
	.out(y3x4_4)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0055196140989170932     ),
	.B1(2*0.0055196140989170932     ),
	.B2(1*0.0055196140989170932     ),
	.A1(-1.7107529570458848       ),
	.A2( 0.73283141344155311      )    
) p4sec4(
	.clk(clk),.en(en),
	.in(y3x4_4),
	.out(y4x5_4)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0055080912957742112     ),
	.B1(2*0.0055080912957742112     ),
	.B2(1*0.0055080912957742112     ),
	.A1(-1.7071815715836276       ),
	.A2( 0.72921393676672441      )    
) p4sec5(
	.clk(clk),.en(en),
	.in(y4x5_4),
	.out(out_4)
);
//part 4 end
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0055004035004604275     ),
	.B1(2*0.0055004035004604275     ),
	.B2(1*0.0055004035004604275     ),
	.A1(-1.7047988110625976       ),
	.A2( 0.72680042506443931      )
) p5sec1 (
	.clk(clk),.en(en),
	.in(out_4),
	.out(y1x2_5)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.0054965578533076086     ),
	.B1(2 *0.0054965578533076086     ),
	.B2(1*0.0054965578533076086     ),
	.A1(-1.7036068885621225       ),
	.A2( 0.72559311997535292      )
) p5sec2 (
	.clk(clk),.en(en),
	.in(y1x2_5),
	.out(out)
);




endmodule 