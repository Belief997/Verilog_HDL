//when put into vivado ,make sure to change the sec1-port-in(in) to in(the_in) 

module my_iir(
	input clk,
	input signed [31:0] in,
	output signed [31:0] out

);
	wire signed [31:0] y1x2, y2x3, y3x4,y4x5,y5x6;
	reg signed [31:0] the_in, sec12, sec23, sec34, sec45, sec56;
	reg [3:0] cnten;
initial begin cnten = 4'b1; the_in = 'b0; sec12 ='b0;sec23 ='b0;sec34 ='b0;sec45 ='b0;sec56 ='b0; end
always @(posedge clk) begin
	if(/*(cnten!= 4'b0)&&*/(cnten!=4'd10))
		cnten <= cnten + 1'b1;
	else if (cnten == 4'd10) begin
		cnten <= 4'd10;
	end 

end

always @(posedge clk) begin
    the_in <= in;
    sec12 <= y1x2;
    sec23 <= y2x3;
    sec34 <= y3x4;
    sec45 <= y4x5;
    sec56 <= y5x6;
end


wire en=(cnten == 4'd10);


////Fs 1K Order 6 Sec3 Elliptic
//IIR_2nd#(
//	.W(32),
//	.FSW(16),
//	.B0(1*0.7961438894),
//	.B1(-1.90032351*0.7961438894),
//	.B2(1*0.7961438894),
//	.A1(-1.885061979),
//	.A2(0.9913290739)
//) sec1 (
//	.clk(clk),.en(en),
//	.in(in),
//	.out(y1x2)
//);
//IIR_2nd#(
//	.W(32),
//	.FSW(16),
//	.B0(1*0.7961438894),
//	.B1(-1.904331803*0.7961438894),
//	.B2(1*0.7961438894),
//	.A1(-1.903072953),
//	.A2(0.9920467138)
//) sec2 (
//	.clk(clk),.en(en),
//	.in(y1x2),
//	.out(y2x3)
//);
//IIR_2nd#(
//	.W(32),
//	.FSW(16),
//	.B0(1*1.526773453),
//	.B1(-1.902347684*1.526773453),
//	.B2(1*1.526773453),
//	.A1(-1.856720924),
//	.A2(0.952031076)
//) sec3 (
//	.clk(clk),.en(en),
//	.in(y2x3),
//	.out(out)
//);
//



////Fs 1k Order 12 Sec 6 Butterworth
//IIR_2nd#(
//	.W(32),
//	.FSW(16),
//	.B0(1*0.99708467737591255),
//	.B1(-1.9023477205076051*0.99708467737591255),
//	.B2(1*0.99708467737591255),
//	.A1(-1.8899259924843124),
//	.A2(0.99409567057051074)
//) sec1 (
//	.clk(clk),.en(en),
//	.in(the_in),
//	.out(y1x2)
//);
//IIR_2nd#(
//	.W(32),
//	.FSW(16),
//	.B0(1*0.99708467737591255),
//	.B1(-1.9023477205076051*0.99708467737591255),
//	.B2(1*0.99708467737591255),
//	.A1(-1.9034616691554653),
//	.A2( 0.99447133786842778)
//) sec2 (
//	.clk(clk),.en(en),
//	.in(sec12),
//	.out(y2x3)
//);
//IIR_2nd#(
//	.W(32),
//	.FSW(16),
//	.B0(1*0.99219872275966292),
//	.B1(-1.9023477205076051*0.99219872275966292),
//	.B2(1*0.99219872275966292),
//	.A1(-1.8822958588945999),
//	.A2( 0.98408618129638525)
//) sec3 (
//	.clk(clk),.en(en),
//	.in(sec23),
//	.out(y3x4)
//);
//IIR_2nd#(
//	.W(32),
//	.FSW(16),
//	.B0(1*0.99219872275966292),
//	.B1(-1.9023477205076051*0.99219872275966292),
//	.B2(1*0.99219872275966292),
//	.A1(-1.8926041104420395),
//	.A2( 0.9848305851346999)    
//) sec4(
//	.clk(clk),.en(en),
//	.in(sec34),
//	.out(y4x5)
//);
//IIR_2nd#(
//	.W(32),
//	.FSW(16),
//	.B0(1*0.98941031509069011),
//	.B1(-1.9023477205076051*0.98941031509069011),
//	.B2(1*0.98941031509069011),
//	.A1(-1.8802666935566985),
//	.A2(  0.97864362026554819)    
//) sec5(
//	.clk(clk),.en(en),
//	.in(sec45),
//	.out(y5x6)
//);
//IIR_2nd#(
//	.W(32),
//	.FSW(16),
//	.B0(1*0.98941031509069011),
//	.B1(-1.9023477205076051*0.98941031509069011),
//	.B2(1*0.98941031509069011),
//	.A1(-1.8841230786926979),
//	.A2( 0.97901393972174411)    
//) sec6(
//	.clk(clk),.en(en),
//	.in(sec56),
//	.out(out)
//);

//////Fs 1K Order 10 Sec5 Elliptic
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.60600827214482633),
	.B1(-1.900087744679229        *0.60600827214482633),
	.B2(1*0.60600827214482633),
	.A1(-1.8891574814809755       ),
	.A2( 0.99655809877856705      )
) sec1 (
	.clk(clk),.en(en),
	.in(the_in),
	.out(y1x2)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.60600827214482633       ),
	.B1(-1.9045578275663106       *0.60600827214482633       ),
	.B2(1*0.60600827214482633       ),
	.A1(-1.9083918557764812       ),
	.A2( 0.99686817128507554      )
) sec2 (
	.clk(clk),.en(en),
	.in(sec12),
	.out(y2x3)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.99044238331821444       ),
	.B1(-1.9009451204244441       *0.99044238331821444       ),
	.B2(1*0.99044238331821444       ),
	.A1(-1.870140143253431        ),
	.A2( 0.98012895245820342      )
) sec3 (
	.clk(clk),.en(en),
	.in(sec23),
	.out(y3x4)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*0.99044238331821444       ),
	.B1(-1.9037309501415742       *0.99044238331821444       ),
	.B2(1*0.99044238331821444       ),
	.A1(-1.8974097046890916       ),
	.A2( 0.98245934724818818      )    
) sec4(
	.clk(clk),.en(en),
	.in(sec34),
	.out(y4x5)
);
IIR_2nd#(
	.W(32),
	.FSW(16),
	.B0(1*2.6024903490653259        ),
	.B1(-1.9023477205076051       *2.6024903490653259        ),
	.B2(1*2.6024903490653259        ),
	.A1(-1.8245736860102928       ),
	.A2( 0.91823362925831475      )    
) sec5(
	.clk(clk),.en(en),
	.in(sec45),
	.out(out)
);



endmodule 
